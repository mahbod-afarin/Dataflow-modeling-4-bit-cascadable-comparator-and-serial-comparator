library verilog;
use verilog.vl_types.all;
entity test_serial_comp is
end test_serial_comp;
