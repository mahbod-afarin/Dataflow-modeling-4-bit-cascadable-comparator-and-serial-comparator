library verilog;
use verilog.vl_types.all;
entity test_comp_6bit is
end test_comp_6bit;
