library verilog;
use verilog.vl_types.all;
entity test_comp_1bit is
end test_comp_1bit;
